module IM(
 	input [31:0] Addr_in,//the value is the address of running instruction 
 	output reg [31:0] Instruction//run instruction
);
	integer i;
	reg [31:0]Instr[199:0];//Creat 200 Instruction address each is 32-bit


always@(Addr_in)begin
	Instruction=Instr[Addr_in/4];//the address of instruction is 4times
end

initial begin
	for(i=0;i<200;i=i+1)begin
		Instr[i]=32'd0;
	end	

	Instr[0]=32'b010100_01000_01001_01000_00000_010101;//add $t0, $t0, $t1
	Instr[1]=32'b010100_01010_01100_01001_00000_010110;//sub $t1, $t2, $t4
	Instr[2]=32'b010100_01101_00000_01100_00001_010111;//srl $t4, $t5, 1
	Instr[3]=32'b010100_01111_00000_01110_00100_011000;//sll $t6, $t7, 4
	Instr[4]=32'b010100_01001_01010_01011_00000_011001;//xor $t3, $t1, $t2
	Instr[5]=32'b010100_01010_01100_01101_00000_011010;//and $t5, $t4, $t2

	Instr[6]=32'b101011_01111_01000_0000000000000010;//sw $t0, 2($t7) 
	Instr[7]=32'b100011_01111_10001_0000000000000010;//lw $s1, 2($t7)
	Instr[8]=32'b100011_01111_10010_0000000000000100;//lw $s2, 4($t7)
	Instr[9]=32'b101011_01010_01000_0000000000000010;//sw $t0, 2($t2)
	Instr[10]=32'b101011_01001_10011_0000000000000100;//sw $s3, 4($t1)
	Instr[11]=32'b001000_10011_10100_0000000001101111;//addi $s4, $s3, 111
	Instr[12]=32'b001000_10101_10110_0000000000011011;//addi $s6, $s5, 27
	Instr[13]=32'b001001_10110_10001_0000000000001001;//subi $s1, $s6, 9
	Instr[14]=32'b001001_10001_10111_0000000000000101;//subi $s7, $s1, 5

	Instr[15]=32'b000100_11000_11001_0000000000000100;//beq $t8, $t9, 4
	Instr[16]=32'b000100_01100_11000_0000000000000001;//beq $t4, $t8, 1
	Instr[17]=32'b000100_10011_10101_0000000000000100;//beq $s3, $s5, 4
	Instr[18]=32'b000100_01100_01101_0000000000000001;//beq $t4, $t5, 1
	Instr[19]=32'b000010_00000000000000000001111101;//j 125
	Instr[20]=32'b000010_00000000000000000000010000;//j 16

	/*Instr[0]=32'b001000_00000_01000_0000000110111100;//addi $t0, $zero, 444
	Instr[1]=32'b001000_00000_01001_0000001000101011;//addi $t1, $zero, 555
	Instr[2]=32'b001000_01000_01000_0000000011011110;//addi $t0, $t0, 222
	Instr[3]=32'b001001_01001_01001_0000000001101111;//subi $t1, $t1, 111
	Instr[4]=32'b010100_01001_01000_01011_00000_011011;//slt $t3, $t1, $t0
	Instr[5]=32'b000100_00000_01011_0000000000000010;//beq $zero, $t3, 2
	Instr[6]=32'b001000_00000_01010_0000001010011010;//addi $t2, $zero, 666
	Instr[7]=32'b000010_00000000000000000000001001;//j 9
	Instr[8]=32'b001000_00000_01010_0000001100001001;//addi $t2, $zero, 777
	Instr[9]=32'b000010_00000000000000000000000000;//j 0*/

end
endmodule
